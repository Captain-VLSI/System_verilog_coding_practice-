//

module traffic_light;
  typedef enum = {red,green, yello} light_e;
  light_e traffic colours;
